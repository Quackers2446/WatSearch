`timescale 1ns/1ps

module low_swing_tx (
    input logic i,
    output logic c
);

assign c = i;

endmodule

