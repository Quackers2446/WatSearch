`timescale 1ns/1ps


module low_swing_rx (
    input logic i,
    output logic o
);

assign o = i;

endmodule
